

module PYTEST(
    input  wire VDD,
    input  wire VSS,
    input  wire vin,
    output wire vout
);

endmodule
